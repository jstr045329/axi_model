package axi_model_pkg;

`include "axi_model.svh"
`include "axi_master_model.svh"
`include "axi_slave_model.svh"

endpackage

